module Control #(
    parameter SIZE = 32,
    parameter ADDR_W = $clog2(SIZE),
    parameter DATA_W = 32,
    parameter MAC_W = 64
) (

);

endmodule