`include "param.hv"

module Control (
    input wire clk
);

endmodule